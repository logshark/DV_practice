import uvm_pkg::*;

module tb;
    initial begin


        uvm_report_info("TEST","hello world");

    end

endmodule